//-------------------------------------------------------------------------
//    Ball.sv                                                            --
//    Viral Mehta                                                        --
//    Spring 2005                                                        --
//                                                                       --
//    Modified by Stephen Kempf 03-01-2006                               --
//                              03-12-2007                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Modified by Po-Han Huang  03-03-2017                               --
//    Spring 2017 Distribution                                           --
//                                                                       --
//    For use with ECE 298 Lab 7                                         --
//    UIUC ECE Department                                                --
//-------------------------------------------------------------------------


module  ball ( input         Reset, 
                             frame_clk,          // The clock indicating a new frame (~60Hz)
                    input logic [15:0] key,
               output [9:0]  BallX, BallY, BallS // Ball coordinates and size
              );
    
    logic [9:0] Ball_X_Pos, Ball_X_Motion, Ball_Y_Pos, Ball_Y_Motion;
    logic [9:0] Ball_X_Pos_in, Ball_X_Motion_in, Ball_Y_Pos_in, Ball_Y_Motion_in;
    logic jump;
     
    parameter [9:0] Ball_X_Center=320;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center=240;  // Center position on the Y axis
    parameter [9:0] Ball_X_Min=0;       // Leftmost point on the X axis
    parameter [9:0] Ball_X_Max=639;     // Rightmost point on the X axis
    parameter [9:0] Ball_Y_Min=0;       // Topmost point on the Y axis
    parameter [9:0] Ball_Y_Max=479;     // Bottommost point on the Y axis
    parameter [9:0] Ball_X_Step=1;      // Step size on the X axis
    parameter [9:0] Ball_Y_Step=1;      // Step size on the Y axis
    parameter [9:0] Ball_Size=4;        // Ball size
    parameter [9:0] jump_limit=100; 
    
    assign BallX = Ball_X_Pos;
    assign BallY = Ball_Y_Pos;
    assign BallS = Ball_Size;
    
    always_ff @ (posedge frame_clk or posedge Reset)
    begin
        if (Reset)
        begin
            Ball_X_Pos <= Ball_X_Center;
            Ball_Y_Pos <= Ball_Y_Center;
            Ball_X_Motion <= 10'd0;
            Ball_Y_Motion <= 10'd0;
        end
        else 
        begin
            Ball_X_Pos <= Ball_X_Pos_in;
            Ball_Y_Pos <= Ball_Y_Pos_in;
            Ball_X_Motion <= Ball_X_Motion_in;
            Ball_Y_Motion <= Ball_Y_Motion_in;
        end
    end
    
    always_comb
    begin
        // By default, keep motion unchanged
        Ball_X_Motion_in = Ball_X_Motion;
        Ball_Y_Motion_in = Ball_Y_Motion;
        
          // W - up = 001A; 
          // D - right = 0007;
          // A - left = 0004;
          // S - down = 0016;
          case (key)
                // up
                16'h001A: begin
                    Ball_Y_Motion_in = (~(Ball_Y_Step) + 1'b1);
                    // prevent diagonal motion
                    Ball_X_Motion_in = 0;
                    if(jump == 0)
                        jump = 1
                end
                // left
                16'h0007: begin
                    Ball_X_Motion_in = Ball_X_Step;
                    // prevent diagonal motion
                    Ball_Y_Motion_in = 0;
                end
                // right
                16'h0004: begin
                    Ball_X_Motion_in = (~(Ball_Y_Step) + 1'b1);
                    // prevent diagonal motion
                    Ball_Y_Motion_in = 0;
                end
                default:
                    Ball_Y_Motion_in = Ball_Y_Step;
          
          endcase
          
          
          
          
        // Be careful when using comparators with "logic" datatype becuase compiler treats 
        //   both sides of the operator UNSIGNED numbers. (unless with further type casting)
        // e.g. Ball_Y_Pos - Ball_Size <= Ball_Y_Min 
        // If Ball_Y_Pos is 0, then Ball_Y_Pos - Ball_Size will not be -4, but rather a large positive number.

        if( Ball_Y_Pos + Ball_Size = Ball_Y_Max ) begin  // Ball is at the bottom edge, stay and set jump to 0
            Ball_Y_Motion_in = 0;
            jump = 0;
        end

        else if ( Ball_X_Pos + Ball_Size = Ball_X_Max) // ball is at right edge, stay
            Ball_X_Motion_in = 0;

        else if ( Ball_X_Pos = Ball_X_Min + Ball_Size ) // ball is at left edge, stay
            Ball_X_Motion_in = 0;

        else begin
            end

        if(jump == 1) begin
            // Haven't hit jump limit yet, keep going up 
            if(Ball_Y_Pos > jump_limit)
                Ball_Y_Motion_in = (~(Ball_Y_Step) - 1'b1)
            else begin
                Ball_Y_Motion_in = (~(Ball_Y_Step) + 1'b1)
            end
        end


          
          
        // Update the ball's position with its motion
        Ball_X_Pos_in = Ball_X_Pos + Ball_X_Motion;
        Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;
        
    /**************************************************************************************
        ATTENTION! Please answer the following quesiton in your lab report! Points will be allocated for the answers!
        Hidden Question #2/2:
          Notice that Ball_Y_Pos is updated using Ball_Y_Motion. 
          Will the new value of Ball_Y_Motion be used when Ball_Y_Pos is updated, or the old? 
          What is the difference between writing
            "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion;" and 
            "Ball_Y_Pos_in = Ball_Y_Pos + Ball_Y_Motion_in;"?
          How will this impact behavior of the ball during a bounce, and how might that interact with a response to a keypress?
          Give an answer in your Post-Lab.
    **************************************************************************************/
        
    end
    
endmodule
